 
module mux_4_1_gatelevel(
input d1,d2,d3,d4,
input s1,s2,
output y
);




endmodule

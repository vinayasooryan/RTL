


module mux_4_1_behavioral_tb;
input i;

    
endmodule

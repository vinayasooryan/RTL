

module mux_2_1_gatelevel(
input d1,d2,
input s,
output reg y
);
wire w1,w2,w3;
and a1(w1,d2,s);
not
and a2(

endmodule
